`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company          : Semicon_Academi
// Engineer         : Jiyun_Han
// 
// Create Date	    : 2025/09/19
// Design Name      : RV32I
// Module Name      : Inst_ROM
// Target Devices   : Basys3
// Tool Versions    : 2020.2
// Description      : Instrucion ROM
//////////////////////////////////////////////////////////////////////////////////

module Inst_ROM(
    input   logic   [31:0]  iRdAddr,

    output  logic   [31:0]  oRdData
    );

    // Reg & Wire - Logic
    logic   [31:0]  rRom[0:63];

    initial
    begin
    //     // Funct7_Rs2_Rs1_Funct3_Rd_Opcode - R_Type (Rd = Rs1 OP Rs2)
    //     rRom[0]     = 32'b0000000_00010_00001_000_00111_0110011;    // add  x7, x1,  x2     (1 + 2 = 3     -> REG[7])
    //     rRom[1]     = 32'b0100000_01000_01001_000_00111_0110011;    // sub  x7, x9,  x8     (9 - 8 = 1     -> REG[7])
    //     rRom[2]     = 32'b0000000_00001_01000_001_00111_0110011;    // sll  x7, x8,  x1     (8 << 1 = 16   -> REG[7]) 
    //     rRom[3]     = 32'b0000000_00001_01000_101_00111_0110011;    // srl  x7, x8,  x1     (8 >> 1 = 4    -> REG[7])
    //     rRom[4]     = 32'b0100000_00010_01010_101_00111_0110011;    // sra  x7, x10, x2     (32'hf0_00_00_00 >>> 2 = 32'hfc_00_00_00 -> REG[7]) 
    //     rRom[5]     = 32'b0000000_01010_01011_010_00111_0110011;    // slt  x7, x11, x10    (32'hff_00_00_00 < 32'hf0_00_00_00 = 0   -> REG[7])
    //     rRom[6]     = 32'b0000000_01011_01010_011_00111_0110011;    // sltu x7, x10, x11    (32'hff_00_00_00 < 32'hf0_00_00_00 = 1   -> REG[7])
    //     rRom[7]     = 32'b0000000_01110_01000_100_00111_0110011;    // xor  x7, x8,  x14    (1000 ^ 1110 = 0110 (6)  -> REG[7]) 
    //     rRom[8]     = 32'b0000000_01110_01000_110_00111_0110011;    // or   x7, x8,  x14    (1000 | 1110 = 1110 (14) -> REG[7])
    //     rRom[9]     = 32'b0000000_01110_01000_111_00111_0110011;    // and  x7, x8,  x14    (1000 & 1110 = 1000 (8)  -> REG[7])

    //     // Imm_Rs2_Rs1_Funct3_Imm_Opcode - S_Type (MEM[Rs1+imm] = Rs2)
    //     rRom[10]    = 32'b0000000_10010_01111_010_00101_0100011;    // sw   x18, 5(x5)      (Store Word 15+5 -> x20 = 32'hdd_dd_dd_dd -> RAM[5])
    //     rRom[11]    = 32'b0000000_10011_10000_001_00100_0100011;    // sh   x19, 4(x5)      (Store Half 16+4 -> x20 = 32'hdd_dd_ee_ee -> RAM[5])
    //     rRom[12]    = 32'b0000000_10011_10000_001_00110_0100011;    // sh   x19, 6(x5)      (Store Half 16+6 -> x22 = 32'hee_ee_ee_ee -> RAM[5])
    //     rRom[13]    = 32'b0000000_10100_10001_000_00011_0100011;    // sb   x20, 3(x5)      (Store Byte 17+3 -> x20 = 32'hee_ee_ee_ff -> RAM[5])
    //     rRom[14]    = 32'b0000000_10100_10001_000_00100_0100011;    // sb   x20, 4(x5)      (Store Byte 17+4 -> x21 = 32'hee_ee_ff_ff -> RAM[5])
    //     rRom[15]    = 32'b0000000_10100_10001_000_00101_0100011;    // sb   x20, 5(x5)      (Store Byte 17+5 -> x22 = 32'hee_ff_ff_ff -> RAM[5])
    //     rRom[16]    = 32'b0000000_10100_10001_000_00110_0100011;    // sb   x20, 6(x5)      (Store Byte 17+6 -> x23 = 32'hff_ff_ff_ff -> RAM[5])

    //     // Imm_Rs1_Funct3_Rd_Opcode - I_Type(L) (Rd = MEM[Rs1 + imm])
    //     rRom[17]    = 32'b000000000000_00100_000_00111_0000011;     // lb   x7, 0(x1)       (Load Byte  32'h00_00_00_21 -> REG[7])
    //     rRom[18]    = 32'b000000000001_00100_000_00111_0000011;     // lb   x7, 1(x1)       (Load Byte  32'h00_00_00_43 -> REG[7])
    //     rRom[19]    = 32'b000000000010_00100_000_00111_0000011;     // lb   x7, 2(x1)       (Load Byte  32'h00_00_00_65 -> REG[7])
    //     rRom[20]    = 32'b000000000011_00100_000_00111_0000011;     // lb   x7, 3(x1)       (Load Byte  32'hff_ff_ff_87 -> REG[7])
    //     rRom[21]    = 32'b000000000011_00101_001_00111_0000011;     // lh   x7, 3(x2)       (Load Byte  32'h00_00_43_22 -> REG[7])
    //     rRom[22]    = 32'b000000000101_00101_001_00111_0000011;     // lh   x7, 5(x2)       (Load Byte  32'hff_ff_87_65 -> REG[7])
    //     rRom[23]    = 32'b000000000110_00110_010_00111_0000011;     // LW   x7, 6(x3)       (Load Byte  32'h87_65_43_23 -> REG[7])
    //     rRom[24]    = 32'b000000000000_00100_100_00111_0000011;     // LBU  x7, 0(x1)       (Load Byte  32'h00_00_00_21 -> REG[7])
    //     rRom[25]    = 32'b000000000001_00100_100_00111_0000011;     // LBU  x7, 1(x1)       (Load Byte  32'h00_00_00_43 -> REG[7])
    //     rRom[26]    = 32'b000000000010_00100_100_00111_0000011;     // LBU  x7, 2(x1)       (Load Byte  32'h00_00_00_65 -> REG[7])
    //     rRom[27]    = 32'b000000000011_00100_100_00111_0000011;     // LBU  x7, 3(x1)       (Load Byte  32'h00_00_00_87 -> REG[7])
    //     rRom[28]    = 32'b000000000011_00101_101_00111_0000011;     // LHU  x7, 3(x2)       (Load Byte  32'h00_00_43_22 -> REG[7])
    //     rRom[29]    = 32'b000000000101_00101_101_00111_0000011;     // LHU  x7, 5(x2)       (Load Byte  32'h00_00_87_65 -> REG[7])

    //     // Imm_Rs1_Funct3_Rd_Opcode - I_Type (Rd = Rs1 OP imm)
    //     rRom[30]    = 32'b000000000010_00001_000_00111_0010011;    // addi  x7, x1,  x2     (1 + 2 = 3     -> REG[7])
    //     rRom[31]    = 32'b000000000001_01000_001_00111_0010011;    // slli  x7, x8,  x1     (8 << 1 = 16   -> REG[7]) 
    //     rRom[32]    = 32'b000000000001_01000_101_00111_0010011;    // srli  x7, x8,  x1     (8 >> 1 = 4    -> REG[7])
    //     rRom[33]    = 32'b010000000010_01010_101_00111_0010011;    // srai  x7, x10, x2     (32'hf0_00_00_00 >>> 2 = 32'hfc_00_00_00 -> REG[7]) 
    //     rRom[34]    = 32'b100000000000_01011_010_00111_0010011;    // slti  x7, x11, x10    (32'hff_00_00_00 < 32'hff_ff_f8_00 = 1   -> REG[7])
    //     rRom[35]    = 32'b100000000000_01010_011_00111_0010011;    // sltiu x7, x10, x11    (32'hff_00_00_00 < 32'h00_00_08_00 = 1   -> REG[7])
    //     rRom[36]    = 32'b000000001110_01000_100_00111_0010011;    // xori  x7, x8,  x14    (1000 ^ 1110 = 0110 (6)  -> REG[7]) 
    //     rRom[37]    = 32'b000000001110_01000_110_00111_0010011;    // ori   x7, x8,  x14    (1000 | 1110 = 1110 (14) -> REG[7])
    //     rRom[38]    = 32'b000000001110_01000_111_00111_0010011;    // andi  x7, x8,  x14    (1000 & 1110 = 1000 (8)  -> REG[7])

    //     // Imm(7)_Rs2_Rs1_Funct3_Imm(5)_Opcode - B_Type (if Rs1 OP Rs2 ? PC : PC + imm)
    //     rRom[39]    = 32'b0000000_00010_00010_000_10000_1100011;    // beq  x2, x2, 16      (2 == 2 Pc+16   -> 43(156 -> 172))
    //     rRom[40]    = 32'b0000000_00001_00010_001_01000_1100011;    // bne  x2, x1, 8       (2 != 1 Pc+8    -> 42(160 -> 168))
    //     rRom[41]    = 32'b0000000_00100_00010_100_10000_1100011;    // blt  x2, x4, 16      (2 <  4 Pc+16   -> 44(164 -> 180))
    //     rRom[42]    = 32'b0000000_00011_00100_101_01000_1100011;    // bge  x4, x3, 8       (4 >= 3 Pc+8    -> 45(168 -> 176))
    //     rRom[43]    = 32'b1111111_00010_00001_110_10101_1100011;    // bltu x1, x2, -12     (1 <  2 Pc-12   -> 40(172 -> 160))
    //     rRom[44]    = 32'b1111111_00010_00011_111_10101_1100011;    // bgeu x3, x2, -12     (3 >= 2 Pc-12   -> 42(176 -> 164))
    //     rRom[45]    = 32'b0000000_00010_00001_000_10000_1100011;    // beq  x1, x2, 16      (1 == 2 Pc+16   -> 46(180 -> 184))
    //     rRom[46]    = 32'b0000000_00010_00010_001_01000_1100011;    // bne  x2, x2, 8       (2 != 2 Pc+8    -> 47(184 -> 188))
    //     rRom[47]    = 32'b0000000_00010_00100_100_10000_1100011;    // blt  x4, x2, 16      (4 <  2 Pc+16   -> 48(188 -> 192))
    //     rRom[48]    = 32'b0000000_00100_00011_101_01000_1100011;    // bge  x3, x4, 8       (3 >= 4 Pc+8    -> 49(192 -> 196))
    //     rRom[49]    = 32'b1111111_00001_00010_110_10101_1100011;    // bltu x2, x1, -12     (2 <  1 Pc-12   -> 50(196 -> 200))
    //     rRom[50]    = 32'b1111111_00011_00010_111_10101_1100011;    // bgeu x2, x3, -12     (2 >= 3 Pc-12   -> 51(200 -> 204))
    //     // 156 -> 172 -> 160 -> 168 -> 176 -> 164 -> 180 -> 184 -> 188 -> 192 -> 196 -> 200 -> 204..

    //     // Imm_Rd_Opcode - U_Type
    //     rRom[51]    = 32'b0000_0000_0000_0001_0100_00111_0110111;   // lui   x7, 0x14       (81920                  -> REG[7])
    //     rRom[52]    = 32'b0000_0000_0000_0001_0100_00111_0010111;   // auipc x7, 0x14       (208 + 81920 = 82128    -> REG[7])

    //     // Imm_Rd_Opcode - JAL (PC += Imm, Rd = PC + 4)
    //     rRom[53]    = 32'b0000_0001_0100_0000_0000_00111_1101111;   // jal  x7, 20          (PC(232) = 212+20,  216 -> REG[7])

    //     // Imm_Rs1_Funct3_Rd_Opcode - JALR (PC = Rs1  + Imm, Rd = PC+4)
    //     rRom[58]    = 32'b000011010000_00100_000_00111_1100111;     // jalr x7  4(x7)       (PC(212) = 4 + 208. 232 -> REG[7] )
    
        $readmemh("code_test1.mem", rRom);
    end
    
    assign  oRdData = rRom[iRdAddr[31:2]];

endmodule